////****\\ Modules to flag events //****\\\\
/*
module Flag (SigFlag, Time, );

//functional I/O's

input [31:0]Time;
input SpikePing;

output [33:0]fList;

//net I/O's

input [7:0]listIndex;

output [7:0]listCount;
endmodule*/
